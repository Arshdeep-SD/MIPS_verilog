`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/16/2020 03:11:42 PM
// Design Name: 
// Module Name: instruction_mem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instruction_mem(
    input [9:0] read_addr,
    output [31:0] data
    );
    
    reg [31:0]rom[255:0];  
    
    initial  
    begin  
                                                        // instruction           alu result in hex       register content       mem content
//        rom[0]  = 32'b00100000000000010000000000000110; // addi r1,r0,#6                 6                    r1=6                   -
//        rom[1]  = 32'b00100000000000100000000000001110; // addi r2,r0,#e                 e                    r2=e                   -
//        rom[2]  = 32'b00100000000000110000000001001110; // addi r3,r0,#4e                4e                   r3=4e                  -
//        rom[3]  = 32'b00100000000001000000000011010010; // addi r4,r0,#d2                d2                   r4=d2                  -
//        rom[4]  = 32'b00100000000001011110000110010101; // addi r5,r0,#e195           ffffe195                r5=ffffe195            -
//        rom[5]  = 32'b00100000000001101111111000010010; // addi r6,r0,#fe12           fffffe12                r6=fffffe12            -
//        rom[6]  = 32'b00000000001001000011100000100000; // add r7,r1,r4                  d8                   r7=d8                  -
//        rom[7]  = 32'b00000000011001010100000000100000; // add r8,r3,r5               ffffe1e3                r8=ffffe1e3            -
//        rom[8]  = 32'b10101100001001110000000000000010; // sw mem[r1+2] <= r7            8                    -                   mem[2]=d8
//        rom[9]  = 32'b10101100100010001111111111111110; // sw mem[r4-2] <= r8            d0                   -                   mem[52]=ffffe1e3
//        rom[10] = 32'b00000000100000100100100000100010; // sub r9,r4,r2                  C4                   r9=c4                  -
//        rom[11] = 32'b00000000001001010101000000100010; // sub r10,r1,r5                1e71                  r10=1e71               -
//        rom[12] = 32'b10101101001010100000000000000000; // sw mem[r9+0] <= r10           c4                   -                   mem[49]=1e71
//        rom[13] = 32'b00000001001001110101100000100101; // or r11,r9,r7                  dc                   r11=dc                 -
//        rom[14] = 32'b00000001000010100110000000100100; // and r12,r8,r10                61                   r12=61                 -
//        rom[15] = 32'b10001100001011010000000000000010; // r13 =mem[r1+2]                8                    r13=d8                 -
//        rom[16] = 32'b10001100100011101111111111111110; // r14 =mem[r4-2]                d0                   r14=ffffe1e3           -
//        rom[17] = 32'b10001101001011110000000000000000; // r15 =mem[r9+0]                c4                   r15=1e71               -
//        rom[18] = 32'b00110001100100000000111101100011; // andi r16,r12,#f63             61                   r16=61                 -
//        rom[19] = 32'b00010000111011010000000000000100; // beq r7,r13,#4                 0                    -                      -              branch to instruction rom[24]     
//        rom[20] = 32'b00000001100010101000100000100111; // nor r17,r12,r10            ffffe18e                r17=ffffe18e           -      
//        rom[21] = 32'b00000001100010101001000000101010; // slt r18,r12,r10               1                    r18=1                  -
//        rom[22] = 32'b11000001100000001001100011000000; // sll r19,r12,#3               308                   r19=308                -
//        rom[23] = 32'b00001000000000000000000000000100; // j #4                          -                    -                      -             jump to instruction rom[28]
//        rom[24] = 32'b11000001100000001010000101000010; // srl r20,r12,#5                3                    r20=3                  -
//        rom[25] = 32'b11000001000000001010100110000011; // sra r21,r8,#6              ffffff87                r21=ffffff87           -
//        rom[26] = 32'b00000000100001011011000000100110; // xor r22,r4,r5              ffffe147                r22=ffffe147           -
//        rom[27] = 32'b00010001010011111111111111111000; // beq r10,r15,#-8                0                   -                      -              branch to instruction rom[20] 
//        rom[28] = 32'b00000000100000011011100000011000; // mult r23,r4,r1                4ec                  r23=4ec                -
//        rom[29] = 32'b00000000111000011100000000011010; // div r24,r7,r1                 24                   r24=24                 -
        
        
        ////////////////////////////////////////////////////// grading
        // load to registers 1 to 10
                                                        // instruction           alu result in hex       register content       mem content
        rom[0] = 32'b10001100000000010000000000000000; // r1  = mem[0]                0                    r1 = 00000001            -
        rom[1] = 32'b10001100000000100000000000000100; // r2  = mem[0]                1                    r2 = 0fd76e10            -
        rom[2] = 32'b10001100000000110000000000001000; // r3  = mem[0]                2                    r3 = 5a00429b            -
        rom[3] = 32'b10001100000001000000000000001100; // r4  = mem[0]                3                    r4 = 14333ffc            -
        rom[4] = 32'b10001100000001010000000000010000; // r5  = mem[0]                4                    r5 = 321fedcb            -
        rom[5] = 32'b10001100000001100000000000010100; // r6  = mem[0]                5                    r6 = 80000000            -
        rom[6] = 32'b10001100000001110000000000011000; // r7  = mem[0]                6                    r7 = 9012fd65            -
        rom[7] = 32'b10001100000010000000000000011100; // r8  = mem[0]                7                    r8 = abc00237            -
        rom[8] = 32'b10001100000010010000000000100000; // r9  = mem[0]                8                    r9 = b54bc031            -
        rom[9] = 32'b10001100000010100000000000100100; // r10 = mem[0]                9                    r10= c187a606            -
        
        // two positive operands
        rom[10] = 32'b00110000011010111111111101100011; // andi r11,r3,#ff63      5a004203                 r11= 5a004203            -
        rom[11] = 32'b00000000001000100110000000100111; // nor  r12,r1,r2         f02891ee                 r12= f02891ee            - 
        rom[12] = 32'b00000000001000100110100000101010; // slt  r13,r1,r2             1                    r13= 1                   -
        rom[13] = 32'b11000000010000000111000011000000; // sll  r14,r2,#3         7ebb7080                 r14= 7ebb7080            -
        rom[14] = 32'b11000000001000000111100101000010; // srl  r15,r1,#5             0                    r15= 0                   -
        rom[15] = 32'b11000000110000001000000110000011; // sra  r16,r6,#6         fe000000                 r16= fe000000            -
        rom[16] = 32'b00000000010000111000100000100110; // xor  r17,r2,r3         55d72c8b                 r17= 55d72c8b            -
        rom[17] = 32'b00000000001000101001000000011000; // mult r17,r1,r2         0fd76e10                 r18= 0fd76e10            -
        rom[18] = 32'b00000000010000011001100000011010; // div  r19,r2,r1         0fd76e10                 r19= 0fd76e10            -
        // store the result in memory
        rom[19] = 32'b10101100000010110000000000101100; // sw mem[r0+11] <= r11      2c                           -                   mem[11]= 5a004203
        rom[20] = 32'b10101100000011000000000000110000; // sw mem[r0+12] <= r12      30                           -                   mem[12]= f02891ee
        rom[21] = 32'b10101100000011010000000000110100; // sw mem[r0+13] <= r13      34                           -                   mem[13]=    1   
        rom[22] = 32'b10101100000011100000000000111000; // sw mem[r0+14] <= r14      38                           -                   mem[14]= 7ebb7080
        rom[23] = 32'b10101100000011110000000000111100; // sw mem[r0+15] <= r15      3c                           -                   mem[15]=    0   
        rom[24] = 32'b10101100000100000000000001000000; // sw mem[r0+16] <= r16      40                          -                   mem[16]= fe000000
        rom[25] = 32'b10101100000100010000000001000100; // sw mem[r0+17] <= r17      44                          -                   mem[17]= 55d72c8b
        rom[26] = 32'b10101100000100100000000001001000; // sw mem[r0+18] <= r18      48                          -                   mem[18]= 0fd76e10
        rom[27] = 32'b10101100000100110000000001001100; // sw mem[r0+19] <= r19      4c                          -                   mem[19]= 0fd76e10
        
        // one positive and one negative operand
        rom[28] = 32'b00110000111010110000111101100011; // andi r11,r7,#f63       00000d61                 r11= 00000d61             -
        rom[29] = 32'b00000000010001110110000000100111; // nor  r12,r2,r7         6028008a                 r12= 6028008a             -
        rom[30] = 32'b00000000010001110110100000101010; // slt  r13,r2,r7             1                    r13=    1                 -
        rom[31] = 32'b11000000111000000111001101000000; // sll  r14,r2,#13        5faca000                 r14= 5faca000             -
        rom[32] = 32'b11000001000000000111100111000010; // srl  r15,r8,#7         01578004                 r15= 01578004             -
        rom[33] = 32'b11000001001000001000000010000011; // sra  r16,r9,#2         ed52f00c                 r16= ed52f00c             -
        rom[34] = 32'b00000000010001111000100000100110; // xor  r17,r2,r7         9fc59375                 r17= 9fc59375             -
        rom[35] = 32'b00000000010001111001000000011000; // mult r17,r2,r7         e4e43c50?                r18= e4e43c50             -
        rom[36] = 32'b00000000111000101001100000011010; // div  r19,r7,r2             9                    r19=    9                 -
        // store the result in memory
        rom[37] = 32'b10101100000010110000000001010000; // sw mem[r0+20] <= r11      50                           -                   mem[20]= 00000d61 
        rom[38] = 32'b10101100000011000000000001010100; // sw mem[r0+21] <= r12      54                           -                   mem[21]= 6028008a 
        rom[39] = 32'b10101100000011010000000001011000; // sw mem[r0+22] <= r13      58                           -                   mem[22]=    1        
        rom[40] = 32'b10101100000011100000000001011100; // sw mem[r0+23] <= r14      5c                           -                   mem[23]= 5faca000 
        rom[41] = 32'b10101100000011110000000001100000; // sw mem[r0+24] <= r15      60                           -                   mem[24]= 01578004 
        rom[42] = 32'b10101100000100000000000001100100; // sw mem[r0+25] <= r16      64                           -                   mem[25]= ed52f00c 
        rom[43] = 32'b10101100000100010000000001101000; // sw mem[r0+26] <= r17      68                           -                   mem[26]= 9fc59375 
        rom[44] = 32'b10101100000100100000000001101100; // sw mem[r0+27] <= r18      6c                           -                   mem[27]= e4e43c50
        rom[45] = 32'b10101100000100110000000001110000; // sw mem[r0+28] <= r19      70                           -                   mem[28]=    9        
        
        // one positive and one negative operand
        rom[46] = 32'b00110001010010111110000100100111; // andi r11,r10,#e127     c187a006                 r11= c187a006             -
        rom[47] = 32'b00000000011010000110000000100111; // nor  r12,r3,r8         043fbd40                 r12= 043fbd40             -
        rom[48] = 32'b00000001000000110110100000101010; // slt  r13,r8,r3             0                    r13=     0                -
        rom[49] = 32'b11000000011000000111010001000000; // sll  r14,r3,#17        85360000                 r14= 85360000             -
        rom[50] = 32'b11000001000000000111110100000010; // srl  r15,r8,#20        00000abc                 r15= 00000abc             -
        rom[51] = 32'b11000001000000001000000001000011; // sra  r16,r8,#1         d5e0011b                 r16= d5e0011b             -
        rom[52] = 32'b00000000011010001000100000100110; // xor  r17,r3,r8         f1c040ac                 r17= f1c040ac             -
        rom[53] = 32'b00000000011010001001000000011000; // mult r17,r3,r8         d3d3854d?                 r18= d3d3854d?             -
        rom[54] = 32'b00000001000000111001100000011010; // div  r19,r8,r3             1                    r19=     1                -
        // store the result in memory
        rom[55] = 32'b10101100000010110000000001110100; // sw mem[r0+29] <= r11      74                           -                   mem[29]= c187a006 
        rom[56] = 32'b10101100000011000000000001111000; // sw mem[r0+30] <= r12      78                           -                   mem[30]= 043fbd40 
        rom[57] = 32'b10101100000011010000000001111100; // sw mem[r0+31] <= r13      7c                           -                   mem[31]=     0       
        rom[58] = 32'b10101100000011100000000010000000; // sw mem[r0+32] <= r14      80                           -                   mem[32]= 85360000 
        rom[59] = 32'b10101100000011110000000010000100; // sw mem[r0+33] <= r15      84                           -                   mem[33]= 00000abc 
        rom[60] = 32'b10101100000100000000000010001000; // sw mem[r0+34] <= r16      88                           -                   mem[34]= d5e0011b 
        rom[61] = 32'b10101100000100010000000010001100; // sw mem[r0+35] <= r17      8c                           -                   mem[35]= f1c040ac 
        rom[62] = 32'b10101100000100100000000010010000; // sw mem[r0+36] <= r18      90                           -                   mem[36]= d3d3854d
        rom[63] = 32'b10101100000100110000000010010100; // sw mem[r0+37] <= r19      94                           -                   mem[37]=     1   

        // two negative operands (not for shift)
        rom[64] = 32'b00110001000010111101000000000010; // andi r11,r8,#d002      abc00002                 r11= abc00002             -
        rom[65] = 32'b00000000111010000110000000100111; // nor  r12,r7,r8         442d0088                 r12= 442d0088             -
        rom[66] = 32'b00000001000001110110100000101010; // slt  r13,r8,r7             0                    r13=     0                -
        rom[67] = 32'b11000000111000000111000111000000; // sll  r14,r7,#7         097eb280                 r14= 097eb280             -
        rom[68] = 32'b11000001001000000111100011000010; // srl  r15,r9,#3         16a97806                 r15= 16a97806             -
        rom[69] = 32'b11000001001000001000000101000011; // sra  r16,r9,#5         fdaa5e01                 r16= fdaa5e01             -
        rom[70] = 32'b00000000111010001000100000100110; // xor  r17,r7,r8         3bd2ff52                 r17= f1c040ac             -
        rom[71] = 32'b00000000111010001001000000011000; // mult r17,r7,r8         9ccf3ab3?                 r18= 9ccf3ab3??             -
        rom[72] = 32'b00000001000001111001100000011010; // div  r19,r8,r7             1                    r19=     1                -
        // store the result in memory
        rom[73] = 32'b10101100000010110000000010011000; // sw mem[r0+38] <= r11      98                           -                   mem[38]= abc00002 
        rom[74] = 32'b10101100000011000000000010011100; // sw mem[r0+39] <= r12      9c                           -                   mem[39]= 442d0088 
        rom[75] = 32'b10101100000011010000000010100000; // sw mem[r0+40] <= r13      a0                           -                   mem[40]=     0       
        rom[76] = 32'b10101100000011100000000010100100; // sw mem[r0+41] <= r14      a4                           -                   mem[41]= 097eb280 
        rom[77] = 32'b10101100000011110000000010101000; // sw mem[r0+42] <= r15      a8                           -                   mem[42]= 16a97806 
        rom[78] = 32'b10101100000100000000000010101100; // sw mem[r0+43] <= r16      ac                           -                   mem[43]= fdaa5e01 
        rom[79] = 32'b10101100000100010000000010110000; // sw mem[r0+44] <= r17      b0                           -                   mem[44]= 3bd2ff52 
        rom[80] = 32'b10101100000100100000000010110100; // sw mem[r0+45] <= r18      b4                           -                   mem[45]= 9ccf3ab3
        rom[81] = 32'b10101100000100110000000010111000; // sw mem[r0+46] <= r19      b8                           -                   mem[46]=     1   

        // zero result or overflow
        rom[82] = 32'b00110001000010110000000000000000; // andi r11,r8,#0         00000000                 r11= 00000000             -
        rom[83] = 32'b00000000110010100110000000100111; // nor  r12,r6,r10        3e7859f9                 r12= 3e7859f9             -
        rom[84] = 32'b00000000110010100110100000101010; // slt  r13,r6,r10            1                    r13=     1                -
        rom[85] = 32'b11000000111000000111011111000000; // sll  r14,r7,#31        80000000                 r14= 80000000             -
        rom[86] = 32'b11000001001000000111111111000010; // srl  r15,r9,#31        00000001                 r15= 00000001             -
        rom[87] = 32'b11000001001000001000011111000011; // sra  r16,r9,#31        ffffffff                 r16= ffffffff             -
        rom[88] = 32'b00000001001010101000100000100110; // xor  r17,r9,r10        74cc6637                 r17= 74cc6637             -
        rom[89] = 32'b00000001001010101001000000011000; // mult r17,r9,r10        a93d4726                 r18= a93d4726??             -
        rom[90] = 32'b00000001001010101001100000011010; // div  r19,r9,r10            0                    r19=     0                -
        // store the result in memory
        rom[91] = 32'b10101100000010110000000010111100; // sw mem[r0+47] <= r11      bc                           -                   mem[47]= 00000000 
        rom[92] = 32'b10101100000011000000000011000000; // sw mem[r0+48] <= r12      c0                           -                   mem[48]= 3e7859f9 
        rom[93] = 32'b10101100000011010000000011000100; // sw mem[r0+49] <= r13      c4                           -                   mem[49]=     1       
        rom[94] = 32'b10101100000011100000000011001000; // sw mem[r0+50] <= r14      c8                           -                   mem[50]= 80000000 
        rom[95] = 32'b10101100000011110000000011001100; // sw mem[r0+51] <= r15      cc                           -                   mem[51]= 00000001 
        rom[96] = 32'b10101100000100000000000011010000; // sw mem[r0+52] <= r16      d0                           -                   mem[52]= ffffffff 
        rom[97] = 32'b10101100000100010000000011010100; // sw mem[r0+53] <= r17      d4                           -                   mem[53]= 74cc6637 
        rom[98] = 32'b10101100000100100000000011011000; // sw mem[r0+54] <= r18      d8                           -                   mem[54]= a93d4726
        rom[99] = 32'b10101100000100110000000011011100; // sw mem[r0+55] <= r19      dc                           -                   mem[55]=     0   


        rom[100] = 32'b00100000001011011111111111111101; // addi r13,r1,#fffd        fffffffe               r13 = fffffffe            -
        rom[101] = 32'b10001100000011100000000000000000; // r14  = mem[0]              0                    r14 = 00000001            -
        rom[102] = 32'b00100000001011111111111111111110; // addi r15,r1,#fffe        ffffffff               r15 = ffffffff            -
         
        
        // branch forward taken
        rom[103] = 32'b00010000001011100000000000000001; // beq r1,r14,#1              0          branch to instruction rom[105]     
        rom[104] = 32'b00000000001000100101000000100000; // add r10,r1,r2         0fd76e11                 r10= 0fd76e11              doesnt run
        rom[105] = 32'b00000000001000111001100000100000; // add r19,r1,r3         5a00429c                 r19= 5a00429c              - 
        rom[106] = 32'b10101100000010100000000011100000; // sw mem[r0+56] <= r10      e0                           -                   mem[56]= c187a606
        
        // branch forward not taken
        rom[107] = 32'b00010000110010100000000000000001; // beq r6,r10,#1         be7859fa        not taken    
        rom[108] = 32'b00000000001001000110000000100000; // add r12,r1,r4         14333ffd                 r12= 14333ffd              
        rom[109] = 32'b00000000001000111001100000100000; // add r19,r1,r3         5a00429c                 r19= 5a00429c              -
        rom[110] = 32'b10101100000011000000000011100100; // sw mem[r0+57] <= r12      e4                           -                   mem[57]= 14333ffd
        
        // branch backward taken
        rom[111] = 32'b00100001101011010000000000000001; // addi r13,r13,#1       ffffffff                                            -  
        rom[112] = 32'b00010001101011111111111111111110; // beq r13,r15,#-2          0            branch to instruction rom[111] 
        // here if the content of r13 = fffffffd then the branch works
        rom[113] = 32'b10101100000011010000000011101000; // sw mem[r0+58] <= r13      e8                           -                   mem[58]= 0
        
        // branch backward not taken
        rom[114] = 32'b00100001110100000000000000000011; // addi r16,r14,#3           4                    r16 = 4                    -       
        rom[115] = 32'b00000010000000011000000000100000; // add r16,r16,r1            5                    r16 = 5                    - 
        rom[116] = 32'b00010000001100001111111111111110; // beq r1,r16,#-2            0            not taken      
//         if the content of r13 = 2 then the branch works
        rom[117] = 32'b10101100000100000000000011101100; // sw mem[r0+59] <= r16      ec                           -                   mem[59]= 5
        
        // branch forward taken
        rom[118] = 32'b00010000001011100000000000000001; // beq r1,r14,#1              0          branch to instruction rom[120]     
        rom[119] = 32'b00000000001000100111100000100000; // add r15,r1,r2         0fd76e11                 r15= 0fd76e11              doesnt run
        rom[120] = 32'b00000000001000111001100000100000; // add r19,r1,r3         5a00429c                 r19= 5a00429c              - 
        rom[121] = 32'b10101100000011110000000011110000; // sw mem[r0+60] <= r15      f0                           -                   mem[60]= ffffffff


        
        //jump forward 
        rom[122] = 32'b00001000000000000000000001111100; // j #7c                    jump to instruction rom[124]          
        rom[123] = 32'b00000000001000100101000000100000; // add r10,r1,r2           0fd76e11                 r10= 0fd76e11       doesnt run         
        rom[124] = 32'b10101100000010100000000011110100; // sw mem[r0+61] <= r10      f4                           -                   mem[61]= c187a606
       
        //jump forward 
        rom[125] = 32'b00001000000000000000000010000000; // j #80                    jump to instruction rom[128]             
        rom[126] = 32'b00000000001000100100100000100000; // add r9,r1,r2          0fd76e11                 r9= 0fd76e11              - 
        rom[127] = 32'b00000000001000100111100000100000; // add r15,r1,r2         0fd76e11                 r15= 0fd76e11        
        rom[128] = 32'b10101100000010010000000011111000; // sw mem[r0+62] <= r9      f8                           -                    mem[62]= b54bc031
        
        //jump forward 
        rom[129] = 32'b00001000000000000000000010000100; // j #84                    jump to instruction rom[132]             
        rom[130] = 32'b00000000001000100100000000100000; // add r8,r1,r2          0fd76e11                 r8= 0fd76e11              - 
        rom[131] = 32'b00000000001000100111100000100000; // add r15,r1,r2         0fd76e11                 r15= 0fd76e11        
        rom[132] = 32'b10101100000010000000000011111100; // sw mem[r0+63] <= r8      fc                           -                    mem[63]= abc00237
        
        //jump forward 
        rom[133] = 32'b00001000000000000000000010001000; // j #88                    jump to instruction rom[132]             
        rom[134] = 32'b00000000001000100011100000100000; // add r7,r1,r2          0fd76e11                 r7= 0fd76e11              - 
        rom[135] = 32'b00000000001000100111100000100000; // add r15,r1,r2         0fd76e11                 r15= 0fd76e11        
        rom[136] = 32'b10101100000001110000000100000000; // sw mem[r0+64] <= r7      100                           -                    mem[64]= 9012fd65
        
        //jump forward 
        rom[137] = 32'b00001000000000000000000010001100; // j #8c                    jump to instruction rom[132]             
        rom[138] = 32'b00000000001000100011000000100000; // add r6,r1,r2          0fd76e11                 r6= 0fd76e11              - 
        rom[139] = 32'b00000000001000100111100000100000; // add r15,r1,r2         0fd76e11                 r15= 0fd76e11        
        rom[140] = 32'b10101100000001100000000100000100; // sw mem[r0+65] <= r6      104                           -                    mem[65]= 80000000
        

        
      end  
      
      assign data = rom[read_addr[9:2]];

endmodule
